module OVERTURE (clk, rst, arch_input_enable, arch_input_value, arch_output_enable, arch_output_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;
  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;

  TC_Switch # (.UUID(64'd3 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_0 (.en(wire_7), .in(arch_input_value), .out(wire_0_6));
  TC_Splitter8 # (.UUID(64'd1677612848903757104 ^ UUID)) Splitter8_1 (.in(wire_1), .out0(wire_28), .out1(wire_5), .out2(wire_40), .out3(wire_23), .out4(wire_17), .out5(wire_6), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd4513427955050900611 ^ UUID)) Decoder3_2 (.dis(wire_26), .sel0(wire_28), .sel1(wire_5), .sel2(wire_40), .out0(wire_8), .out1(wire_21), .out2(wire_32), .out3(wire_22), .out4(wire_38), .out5(wire_31), .out6(wire_19), .out7());
  TC_Decoder3 # (.UUID(64'd3886037073670587034 ^ UUID)) Decoder3_3 (.dis(wire_26), .sel0(wire_23), .sel1(wire_17), .sel2(wire_6), .out0(wire_10), .out1(wire_24), .out2(wire_18), .out3(wire_14), .out4(wire_12), .out5(wire_33), .out6(wire_7), .out7());
  TC_IOSwitch # (.UUID(64'd4 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_4 (.in(wire_0), .en(wire_19), .out(arch_output_value));
  TC_Switch # (.UUID(64'd1031995853711794913 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_16), .in(wire_27), .out(wire_37_0));
  TC_Not # (.UUID(64'd4158910752250590214 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_16), .out(wire_34));
  TC_Switch # (.UUID(64'd4099835737832785551 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_34), .in(wire_0), .out(wire_37_1));
  TC_Xor # (.UUID(64'd3040775265495990141 ^ UUID), .BIT_WIDTH(64'd1)) Xor_8 (.in0(wire_22), .in1(wire_16), .out(wire_20));
  TC_Counter # (.UUID(64'd92340409037022771 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_9 (.clk(clk), .rst(rst), .save(wire_13), .in(wire_9), .out(wire_3));
  TC_Switch # (.UUID(64'd2128825035222160525 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_41), .in(wire_0), .out(wire_11_1));
  TC_Switch # (.UUID(64'd1154064313276925863 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_4), .in(wire_1), .out(wire_11_0));
  TC_Switch # (.UUID(64'd4048984116695642554 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_15), .in(wire_1), .out(wire_25));
  TC_Switch # (.UUID(64'd3052318132109565257 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_13), .in(wire_39), .out(wire_9));
  TC_Not # (.UUID(64'd4481080336099558156 ^ UUID), .BIT_WIDTH(64'd1)) Not_14 (.in(wire_29), .out(wire_26));
  TC_Not # (.UUID(64'd1679235009118185088 ^ UUID), .BIT_WIDTH(64'd1)) Not_15 (.in(wire_4), .out(wire_41));
  TC_Or # (.UUID(64'd4017470350233035878 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_8), .in1(wire_4), .out(wire_36));
  TC_Program8_1 # (.UUID(64'd5 ^ UUID), .DEFAULT_FILE_NAME("Program8_1_5.w8.bin"), .ARG_SIG("Program8_1_5=%s")) Program8_1_17 (.clk(clk), .rst(rst), .address(wire_3), .out(wire_1));
  DEC # (.UUID(64'd3005803602252776583 ^ UUID)) DEC_18 (.clk(clk), .rst(rst), .OPCODE(wire_1), .IMMEDIATE(wire_4), .CALCULATION(wire_16), .COPY(wire_29), .CONDITION(wire_15));
  ALU # (.UUID(64'd1867860043825594088 ^ UUID)) ALU_19 (.clk(clk), .rst(rst), .Instruction(wire_1), .Input_1(wire_30), .Input_2(wire_2), .Output(wire_27));
  COND # (.UUID(64'd3713771086149463027 ^ UUID)) COND_20 (.clk(clk), .rst(rst), .Condition(wire_25), .Input(wire_35), .Result(wire_13));
  RegisterPlus # (.UUID(64'd100000 ^ UUID)) RegisterPlus_21 (.clk(clk), .rst(rst), .Load(wire_10), .Save_value(wire_11), .Save(wire_36), .Always_output(wire_39), .Output(wire_0_5));
  RegisterPlus # (.UUID(64'd110000 ^ UUID)) RegisterPlus_22 (.clk(clk), .rst(rst), .Load(wire_24), .Save_value(wire_0), .Save(wire_21), .Always_output(wire_30), .Output(wire_0_4));
  RegisterPlus # (.UUID(64'd120000 ^ UUID)) RegisterPlus_23 (.clk(clk), .rst(rst), .Load(wire_18), .Save_value(wire_0), .Save(wire_32), .Always_output(wire_2), .Output(wire_0_3));
  RegisterPlus # (.UUID(64'd140000 ^ UUID)) RegisterPlus_24 (.clk(clk), .rst(rst), .Load(wire_12), .Save_value(wire_0), .Save(wire_38), .Always_output(), .Output(wire_0_0));
  RegisterPlus # (.UUID(64'd150000 ^ UUID)) RegisterPlus_25 (.clk(clk), .rst(rst), .Load(wire_33), .Save_value(wire_0), .Save(wire_31), .Always_output(), .Output(wire_0_1));
  RegisterPlus # (.UUID(64'd1161571428188987910 ^ UUID)) RegisterPlus_26 (.clk(clk), .rst(rst), .Load(wire_14), .Save_value(wire_37), .Save(wire_20), .Always_output(wire_35), .Output(wire_0_2));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  wire [7:0] wire_0_4;
  wire [7:0] wire_0_5;
  wire [7:0] wire_0_6;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign arch_input_enable = wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_11_0;
  wire [7:0] wire_11_1;
  assign wire_11 = wire_11_0|wire_11_1;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  assign arch_output_enable = wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_37_0;
  wire [7:0] wire_37_1;
  assign wire_37 = wire_37_0|wire_37_1;
  wire [0:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;

endmodule
